module NOT_G(A,B);
input A;
output B;
assign B=~A;


endmodule